`timescale 1ns / 1ps

module genRandNum(
    input clk
);

always @(posedge clk)
    